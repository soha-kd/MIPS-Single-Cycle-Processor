`timescale 1ns/1ns
module Mux32bit(input [31:0]a, b, input s, output [31:0] w);
	assign w = s == 1'b0 ? a : b;
endmodule
